
module MIPSMonitor (
	source,
	probe);	

	output	[0:0]	source;
	input	[510:0]	probe;
endmodule
